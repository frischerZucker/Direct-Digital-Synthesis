-- Algorithmische Ebense -----------------------------------------------------------------------------------
architecture algorithmisch of dds is

signal f_ref : std_ulogic;					-- Referenzfrequenz mit 48.828 kHz -> Takt f�r Phasenakkumulator
signal phase : integer range 0 to 4095;		-- aktuelle Phase -> Index f�r Koeffiziententabelle
-- Koeffizienten der Funktion
signal coef_table : coef_table_t := (0=>511,1=>512,2=>513,3=>513,4=>514,5=>515,6=>516,7=>516,8=>517,9=>518,10=>519,11=>520,12=>520,13=>521,14=>522,15=>523,16=>524,17=>524,18=>525,19=>526,20=>527,21=>527,22=>528,23=>529,24=>530,25=>531,26=>531,27=>532,28=>533,29=>534,30=>535,31=>535,32=>536,33=>537,34=>538,35=>538,36=>539,37=>540,38=>541,39=>542,40=>542,41=>543,42=>544,43=>545,44=>545,45=>546,46=>547,47=>548,48=>549,49=>549,50=>550,51=>551,52=>552,53=>553,54=>553,55=>554,56=>555,57=>556,58=>556,59=>557,60=>558,61=>559,62=>560,63=>560,64=>561,65=>562,66=>563,67=>563,68=>564,69=>565,70=>566,71=>567,72=>567,73=>568,74=>569,75=>570,76=>570,77=>571,78=>572,79=>573,80=>574,81=>574,82=>575,83=>576,84=>577,85=>578,86=>578,87=>579,88=>580,89=>581,90=>581,91=>582,92=>583,93=>584,94=>585,95=>585,96=>586,97=>587,98=>588,99=>588,100=>589,101=>590,102=>591,103=>591,104=>592,105=>593,106=>594,107=>595,108=>595,109=>596,110=>597,111=>598,112=>598,113=>599,114=>600,115=>601,116=>602,117=>602,118=>603,119=>604,120=>605,121=>605,122=>606,123=>607,124=>608,125=>608,126=>609,127=>610,128=>611,129=>612,130=>612,131=>613,132=>614,133=>615,134=>615,135=>616,136=>617,137=>618,138=>618,139=>619,140=>620,141=>621,142=>622,143=>622,144=>623,145=>624,146=>625,147=>625,148=>626,149=>627,150=>628,151=>628,152=>629,153=>630,154=>631,155=>631,156=>632,157=>633,158=>634,159=>635,160=>635,161=>636,162=>637,163=>638,164=>638,165=>639,166=>640,167=>641,168=>641,169=>642,170=>643,171=>644,172=>644,173=>645,174=>646,175=>647,176=>647,177=>648,178=>649,179=>650,180=>650,181=>651,182=>652,183=>653,184=>653,185=>654,186=>655,187=>656,188=>656,189=>657,190=>658,191=>659,192=>659,193=>660,194=>661,195=>662,196=>662,197=>663,198=>664,199=>665,200=>665,201=>666,202=>667,203=>668,204=>668,205=>669,206=>670,207=>671,208=>671,209=>672,210=>673,211=>674,212=>674,213=>675,214=>676,215=>677,216=>677,217=>678,218=>679,219=>680,220=>680,221=>681,222=>682,223=>683,224=>683,225=>684,226=>685,227=>686,228=>686,229=>687,230=>688,231=>688,232=>689,233=>690,234=>691,235=>691,236=>692,237=>693,238=>694,239=>694,240=>695,241=>696,242=>697,243=>697,244=>698,245=>699,246=>699,247=>700,248=>701,249=>702,250=>702,251=>703,252=>704,253=>705,254=>705,255=>706,256=>707,257=>707,258=>708,259=>709,260=>710,261=>710,262=>711,263=>712,264=>713,265=>713,266=>714,267=>715,268=>715,269=>716,270=>717,271=>718,272=>718,273=>719,274=>720,275=>720,276=>721,277=>722,278=>723,279=>723,280=>724,281=>725,282=>725,283=>726,284=>727,285=>728,286=>728,287=>729,288=>730,289=>730,290=>731,291=>732,292=>733,293=>733,294=>734,295=>735,296=>735,297=>736,298=>737,299=>737,300=>738,301=>739,302=>740,303=>740,304=>741,305=>742,306=>742,307=>743,308=>744,309=>744,310=>745,311=>746,312=>747,313=>747,314=>748,315=>749,316=>749,317=>750,318=>751,319=>751,320=>752,321=>753,322=>754,323=>754,324=>755,325=>756,326=>756,327=>757,328=>758,329=>758,330=>759,331=>760,332=>760,333=>761,334=>762,335=>762,336=>763,337=>764,338=>764,339=>765,340=>766,341=>767,342=>767,343=>768,344=>769,345=>769,346=>770,347=>771,348=>771,349=>772,350=>773,351=>773,352=>774,353=>775,354=>775,355=>776,356=>777,357=>777,358=>778,359=>779,360=>779,361=>780,362=>781,363=>781,364=>782,365=>783,366=>783,367=>784,368=>785,369=>785,370=>786,371=>787,372=>787,373=>788,374=>789,375=>789,376=>790,377=>791,378=>791,379=>792,380=>793,381=>793,382=>794,383=>795,384=>795,385=>796,386=>796,387=>797,388=>798,389=>798,390=>799,391=>800,392=>800,393=>801,394=>802,395=>802,396=>803,397=>804,398=>804,399=>805,400=>806,401=>806,402=>807,403=>807,404=>808,405=>809,406=>809,407=>810,408=>811,409=>811,410=>812,411=>813,412=>813,413=>814,414=>814,415=>815,416=>816,417=>816,418=>817,419=>818,420=>818,421=>819,422=>819,423=>820,424=>821,425=>821,426=>822,427=>823,428=>823,429=>824,430=>824,431=>825,432=>826,433=>826,434=>827,435=>828,436=>828,437=>829,438=>829,439=>830,440=>831,441=>831,442=>832,443=>832,444=>833,445=>834,446=>834,447=>835,448=>835,449=>836,450=>837,451=>837,452=>838,453=>839,454=>839,455=>840,456=>840,457=>841,458=>842,459=>842,460=>843,461=>843,462=>844,463=>845,464=>845,465=>846,466=>846,467=>847,468=>847,469=>848,470=>849,471=>849,472=>850,473=>850,474=>851,475=>852,476=>852,477=>853,478=>853,479=>854,480=>855,481=>855,482=>856,483=>856,484=>857,485=>857,486=>858,487=>859,488=>859,489=>860,490=>860,491=>861,492=>861,493=>862,494=>863,495=>863,496=>864,497=>864,498=>865,499=>865,500=>866,501=>867,502=>867,503=>868,504=>868,505=>869,506=>869,507=>870,508=>870,509=>871,510=>872,511=>872,512=>873,513=>873,514=>874,515=>874,516=>875,517=>875,518=>876,519=>877,520=>877,521=>878,522=>878,523=>879,524=>879,525=>880,526=>880,527=>881,528=>881,529=>882,530=>883,531=>883,532=>884,533=>884,534=>885,535=>885,536=>886,537=>886,538=>887,539=>887,540=>888,541=>888,542=>889,543=>889,544=>890,545=>891,546=>891,547=>892,548=>892,549=>893,550=>893,551=>894,552=>894,553=>895,554=>895,555=>896,556=>896,557=>897,558=>897,559=>898,560=>898,561=>899,562=>899,563=>900,564=>900,565=>901,566=>901,567=>902,568=>902,569=>903,570=>903,571=>904,572=>904,573=>905,574=>905,575=>906,576=>906,577=>907,578=>907,579=>908,580=>908,581=>909,582=>909,583=>910,584=>910,585=>911,586=>911,587=>912,588=>912,589=>913,590=>913,591=>914,592=>914,593=>915,594=>915,595=>916,596=>916,597=>917,598=>917,599=>918,600=>918,601=>919,602=>919,603=>919,604=>920,605=>920,606=>921,607=>921,608=>922,609=>922,610=>923,611=>923,612=>924,613=>924,614=>925,615=>925,616=>926,617=>926,618=>926,619=>927,620=>927,621=>928,622=>928,623=>929,624=>929,625=>930,626=>930,627=>931,628=>931,629=>931,630=>932,631=>932,632=>933,633=>933,634=>934,635=>934,636=>935,637=>935,638=>935,639=>936,640=>936,641=>937,642=>937,643=>938,644=>938,645=>938,646=>939,647=>939,648=>940,649=>940,650=>941,651=>941,652=>941,653=>942,654=>942,655=>943,656=>943,657=>944,658=>944,659=>944,660=>945,661=>945,662=>946,663=>946,664=>946,665=>947,666=>947,667=>948,668=>948,669=>949,670=>949,671=>949,672=>950,673=>950,674=>951,675=>951,676=>951,677=>952,678=>952,679=>953,680=>953,681=>953,682=>954,683=>954,684=>954,685=>955,686=>955,687=>956,688=>956,689=>956,690=>957,691=>957,692=>958,693=>958,694=>958,695=>959,696=>959,697=>959,698=>960,699=>960,700=>961,701=>961,702=>961,703=>962,704=>962,705=>962,706=>963,707=>963,708=>964,709=>964,710=>964,711=>965,712=>965,713=>965,714=>966,715=>966,716=>966,717=>967,718=>967,719=>968,720=>968,721=>968,722=>969,723=>969,724=>969,725=>970,726=>970,727=>970,728=>971,729=>971,730=>971,731=>972,732=>972,733=>972,734=>973,735=>973,736=>973,737=>974,738=>974,739=>974,740=>975,741=>975,742=>975,743=>976,744=>976,745=>976,746=>977,747=>977,748=>977,749=>978,750=>978,751=>978,752=>979,753=>979,754=>979,755=>980,756=>980,757=>980,758=>981,759=>981,760=>981,761=>981,762=>982,763=>982,764=>982,765=>983,766=>983,767=>983,768=>984,769=>984,770=>984,771=>984,772=>985,773=>985,774=>985,775=>986,776=>986,777=>986,778=>987,779=>987,780=>987,781=>987,782=>988,783=>988,784=>988,785=>989,786=>989,787=>989,788=>989,789=>990,790=>990,791=>990,792=>990,793=>991,794=>991,795=>991,796=>992,797=>992,798=>992,799=>992,800=>993,801=>993,802=>993,803=>993,804=>994,805=>994,806=>994,807=>994,808=>995,809=>995,810=>995,811=>995,812=>996,813=>996,814=>996,815=>996,816=>997,817=>997,818=>997,819=>997,820=>998,821=>998,822=>998,823=>998,824=>999,825=>999,826=>999,827=>999,828=>1000,829=>1000,830=>1000,831=>1000,832=>1000,833=>1001,834=>1001,835=>1001,836=>1001,837=>1002,838=>1002,839=>1002,840=>1002,841=>1002,842=>1003,843=>1003,844=>1003,845=>1003,846=>1004,847=>1004,848=>1004,849=>1004,850=>1004,851=>1005,852=>1005,853=>1005,854=>1005,855=>1005,856=>1006,857=>1006,858=>1006,859=>1006,860=>1006,861=>1007,862=>1007,863=>1007,864=>1007,865=>1007,866=>1008,867=>1008,868=>1008,869=>1008,870=>1008,871=>1008,872=>1009,873=>1009,874=>1009,875=>1009,876=>1009,877=>1010,878=>1010,879=>1010,880=>1010,881=>1010,882=>1010,883=>1011,884=>1011,885=>1011,886=>1011,887=>1011,888=>1011,889=>1012,890=>1012,891=>1012,892=>1012,893=>1012,894=>1012,895=>1013,896=>1013,897=>1013,898=>1013,899=>1013,900=>1013,901=>1013,902=>1014,903=>1014,904=>1014,905=>1014,906=>1014,907=>1014,908=>1014,909=>1015,910=>1015,911=>1015,912=>1015,913=>1015,914=>1015,915=>1015,916=>1015,917=>1016,918=>1016,919=>1016,920=>1016,921=>1016,922=>1016,923=>1016,924=>1016,925=>1017,926=>1017,927=>1017,928=>1017,929=>1017,930=>1017,931=>1017,932=>1017,933=>1018,934=>1018,935=>1018,936=>1018,937=>1018,938=>1018,939=>1018,940=>1018,941=>1018,942=>1018,943=>1019,944=>1019,945=>1019,946=>1019,947=>1019,948=>1019,949=>1019,950=>1019,951=>1019,952=>1019,953=>1019,954=>1020,955=>1020,956=>1020,957=>1020,958=>1020,959=>1020,960=>1020,961=>1020,962=>1020,963=>1020,964=>1020,965=>1020,966=>1020,967=>1021,968=>1021,969=>1021,970=>1021,971=>1021,972=>1021,973=>1021,974=>1021,975=>1021,976=>1021,977=>1021,978=>1021,979=>1021,980=>1021,981=>1021,982=>1021,983=>1021,984=>1022,985=>1022,986=>1022,987=>1022,988=>1022,989=>1022,990=>1022,991=>1022,992=>1022,993=>1022,994=>1022,995=>1022,996=>1022,997=>1022,998=>1022,999=>1022,1000=>1022,1001=>1022,1002=>1022,1003=>1022,1004=>1022,1005=>1022,1006=>1022,1007=>1022,1008=>1022,1009=>1022,1010=>1022,1011=>1022,1012=>1022,1013=>1022,1014=>1022,1015=>1022,1016=>1022,1017=>1022,1018=>1022,1019=>1022,1020=>1022,1021=>1022,1022=>1022,1023=>1022,1024=>1023,1025=>1022,1026=>1022,1027=>1022,1028=>1022,1029=>1022,1030=>1022,1031=>1022,1032=>1022,1033=>1022,1034=>1022,1035=>1022,1036=>1022,1037=>1022,1038=>1022,1039=>1022,1040=>1022,1041=>1022,1042=>1022,1043=>1022,1044=>1022,1045=>1022,1046=>1022,1047=>1022,1048=>1022,1049=>1022,1050=>1022,1051=>1022,1052=>1022,1053=>1022,1054=>1022,1055=>1022,1056=>1022,1057=>1022,1058=>1022,1059=>1022,1060=>1022,1061=>1022,1062=>1022,1063=>1022,1064=>1022,1065=>1021,1066=>1021,1067=>1021,1068=>1021,1069=>1021,1070=>1021,1071=>1021,1072=>1021,1073=>1021,1074=>1021,1075=>1021,1076=>1021,1077=>1021,1078=>1021,1079=>1021,1080=>1021,1081=>1021,1082=>1020,1083=>1020,1084=>1020,1085=>1020,1086=>1020,1087=>1020,1088=>1020,1089=>1020,1090=>1020,1091=>1020,1092=>1020,1093=>1020,1094=>1020,1095=>1019,1096=>1019,1097=>1019,1098=>1019,1099=>1019,1100=>1019,1101=>1019,1102=>1019,1103=>1019,1104=>1019,1105=>1019,1106=>1018,1107=>1018,1108=>1018,1109=>1018,1110=>1018,1111=>1018,1112=>1018,1113=>1018,1114=>1018,1115=>1018,1116=>1017,1117=>1017,1118=>1017,1119=>1017,1120=>1017,1121=>1017,1122=>1017,1123=>1017,1124=>1016,1125=>1016,1126=>1016,1127=>1016,1128=>1016,1129=>1016,1130=>1016,1131=>1016,1132=>1015,1133=>1015,1134=>1015,1135=>1015,1136=>1015,1137=>1015,1138=>1015,1139=>1015,1140=>1014,1141=>1014,1142=>1014,1143=>1014,1144=>1014,1145=>1014,1146=>1014,1147=>1013,1148=>1013,1149=>1013,1150=>1013,1151=>1013,1152=>1013,1153=>1013,1154=>1012,1155=>1012,1156=>1012,1157=>1012,1158=>1012,1159=>1012,1160=>1011,1161=>1011,1162=>1011,1163=>1011,1164=>1011,1165=>1011,1166=>1010,1167=>1010,1168=>1010,1169=>1010,1170=>1010,1171=>1010,1172=>1009,1173=>1009,1174=>1009,1175=>1009,1176=>1009,1177=>1008,1178=>1008,1179=>1008,1180=>1008,1181=>1008,1182=>1008,1183=>1007,1184=>1007,1185=>1007,1186=>1007,1187=>1007,1188=>1006,1189=>1006,1190=>1006,1191=>1006,1192=>1006,1193=>1005,1194=>1005,1195=>1005,1196=>1005,1197=>1005,1198=>1004,1199=>1004,1200=>1004,1201=>1004,1202=>1004,1203=>1003,1204=>1003,1205=>1003,1206=>1003,1207=>1002,1208=>1002,1209=>1002,1210=>1002,1211=>1002,1212=>1001,1213=>1001,1214=>1001,1215=>1001,1216=>1000,1217=>1000,1218=>1000,1219=>1000,1220=>1000,1221=>999,1222=>999,1223=>999,1224=>999,1225=>998,1226=>998,1227=>998,1228=>998,1229=>997,1230=>997,1231=>997,1232=>997,1233=>996,1234=>996,1235=>996,1236=>996,1237=>995,1238=>995,1239=>995,1240=>995,1241=>994,1242=>994,1243=>994,1244=>994,1245=>993,1246=>993,1247=>993,1248=>993,1249=>992,1250=>992,1251=>992,1252=>992,1253=>991,1254=>991,1255=>991,1256=>990,1257=>990,1258=>990,1259=>990,1260=>989,1261=>989,1262=>989,1263=>989,1264=>988,1265=>988,1266=>988,1267=>987,1268=>987,1269=>987,1270=>987,1271=>986,1272=>986,1273=>986,1274=>985,1275=>985,1276=>985,1277=>984,1278=>984,1279=>984,1280=>984,1281=>983,1282=>983,1283=>983,1284=>982,1285=>982,1286=>982,1287=>981,1288=>981,1289=>981,1290=>981,1291=>980,1292=>980,1293=>980,1294=>979,1295=>979,1296=>979,1297=>978,1298=>978,1299=>978,1300=>977,1301=>977,1302=>977,1303=>976,1304=>976,1305=>976,1306=>975,1307=>975,1308=>975,1309=>974,1310=>974,1311=>974,1312=>973,1313=>973,1314=>973,1315=>972,1316=>972,1317=>972,1318=>971,1319=>971,1320=>971,1321=>970,1322=>970,1323=>970,1324=>969,1325=>969,1326=>969,1327=>968,1328=>968,1329=>968,1330=>967,1331=>967,1332=>966,1333=>966,1334=>966,1335=>965,1336=>965,1337=>965,1338=>964,1339=>964,1340=>964,1341=>963,1342=>963,1343=>962,1344=>962,1345=>962,1346=>961,1347=>961,1348=>961,1349=>960,1350=>960,1351=>959,1352=>959,1353=>959,1354=>958,1355=>958,1356=>958,1357=>957,1358=>957,1359=>956,1360=>956,1361=>956,1362=>955,1363=>955,1364=>954,1365=>954,1366=>954,1367=>953,1368=>953,1369=>953,1370=>952,1371=>952,1372=>951,1373=>951,1374=>951,1375=>950,1376=>950,1377=>949,1378=>949,1379=>949,1380=>948,1381=>948,1382=>947,1383=>947,1384=>946,1385=>946,1386=>946,1387=>945,1388=>945,1389=>944,1390=>944,1391=>944,1392=>943,1393=>943,1394=>942,1395=>942,1396=>941,1397=>941,1398=>941,1399=>940,1400=>940,1401=>939,1402=>939,1403=>938,1404=>938,1405=>938,1406=>937,1407=>937,1408=>936,1409=>936,1410=>935,1411=>935,1412=>935,1413=>934,1414=>934,1415=>933,1416=>933,1417=>932,1418=>932,1419=>931,1420=>931,1421=>931,1422=>930,1423=>930,1424=>929,1425=>929,1426=>928,1427=>928,1428=>927,1429=>927,1430=>926,1431=>926,1432=>926,1433=>925,1434=>925,1435=>924,1436=>924,1437=>923,1438=>923,1439=>922,1440=>922,1441=>921,1442=>921,1443=>920,1444=>920,1445=>919,1446=>919,1447=>919,1448=>918,1449=>918,1450=>917,1451=>917,1452=>916,1453=>916,1454=>915,1455=>915,1456=>914,1457=>914,1458=>913,1459=>913,1460=>912,1461=>912,1462=>911,1463=>911,1464=>910,1465=>910,1466=>909,1467=>909,1468=>908,1469=>908,1470=>907,1471=>907,1472=>906,1473=>906,1474=>905,1475=>905,1476=>904,1477=>904,1478=>903,1479=>903,1480=>902,1481=>902,1482=>901,1483=>901,1484=>900,1485=>900,1486=>899,1487=>899,1488=>898,1489=>898,1490=>897,1491=>897,1492=>896,1493=>896,1494=>895,1495=>895,1496=>894,1497=>894,1498=>893,1499=>893,1500=>892,1501=>892,1502=>891,1503=>891,1504=>890,1505=>889,1506=>889,1507=>888,1508=>888,1509=>887,1510=>887,1511=>886,1512=>886,1513=>885,1514=>885,1515=>884,1516=>884,1517=>883,1518=>883,1519=>882,1520=>881,1521=>881,1522=>880,1523=>880,1524=>879,1525=>879,1526=>878,1527=>878,1528=>877,1529=>877,1530=>876,1531=>875,1532=>875,1533=>874,1534=>874,1535=>873,1536=>873,1537=>872,1538=>872,1539=>871,1540=>870,1541=>870,1542=>869,1543=>869,1544=>868,1545=>868,1546=>867,1547=>867,1548=>866,1549=>865,1550=>865,1551=>864,1552=>864,1553=>863,1554=>863,1555=>862,1556=>861,1557=>861,1558=>860,1559=>860,1560=>859,1561=>859,1562=>858,1563=>857,1564=>857,1565=>856,1566=>856,1567=>855,1568=>855,1569=>854,1570=>853,1571=>853,1572=>852,1573=>852,1574=>851,1575=>850,1576=>850,1577=>849,1578=>849,1579=>848,1580=>847,1581=>847,1582=>846,1583=>846,1584=>845,1585=>845,1586=>844,1587=>843,1588=>843,1589=>842,1590=>842,1591=>841,1592=>840,1593=>840,1594=>839,1595=>839,1596=>838,1597=>837,1598=>837,1599=>836,1600=>835,1601=>835,1602=>834,1603=>834,1604=>833,1605=>832,1606=>832,1607=>831,1608=>831,1609=>830,1610=>829,1611=>829,1612=>828,1613=>828,1614=>827,1615=>826,1616=>826,1617=>825,1618=>824,1619=>824,1620=>823,1621=>823,1622=>822,1623=>821,1624=>821,1625=>820,1626=>819,1627=>819,1628=>818,1629=>818,1630=>817,1631=>816,1632=>816,1633=>815,1634=>814,1635=>814,1636=>813,1637=>813,1638=>812,1639=>811,1640=>811,1641=>810,1642=>809,1643=>809,1644=>808,1645=>807,1646=>807,1647=>806,1648=>806,1649=>805,1650=>804,1651=>804,1652=>803,1653=>802,1654=>802,1655=>801,1656=>800,1657=>800,1658=>799,1659=>798,1660=>798,1661=>797,1662=>796,1663=>796,1664=>795,1665=>795,1666=>794,1667=>793,1668=>793,1669=>792,1670=>791,1671=>791,1672=>790,1673=>789,1674=>789,1675=>788,1676=>787,1677=>787,1678=>786,1679=>785,1680=>785,1681=>784,1682=>783,1683=>783,1684=>782,1685=>781,1686=>781,1687=>780,1688=>779,1689=>779,1690=>778,1691=>777,1692=>777,1693=>776,1694=>775,1695=>775,1696=>774,1697=>773,1698=>773,1699=>772,1700=>771,1701=>771,1702=>770,1703=>769,1704=>769,1705=>768,1706=>767,1707=>767,1708=>766,1709=>765,1710=>764,1711=>764,1712=>763,1713=>762,1714=>762,1715=>761,1716=>760,1717=>760,1718=>759,1719=>758,1720=>758,1721=>757,1722=>756,1723=>756,1724=>755,1725=>754,1726=>754,1727=>753,1728=>752,1729=>751,1730=>751,1731=>750,1732=>749,1733=>749,1734=>748,1735=>747,1736=>747,1737=>746,1738=>745,1739=>744,1740=>744,1741=>743,1742=>742,1743=>742,1744=>741,1745=>740,1746=>740,1747=>739,1748=>738,1749=>737,1750=>737,1751=>736,1752=>735,1753=>735,1754=>734,1755=>733,1756=>733,1757=>732,1758=>731,1759=>730,1760=>730,1761=>729,1762=>728,1763=>728,1764=>727,1765=>726,1766=>725,1767=>725,1768=>724,1769=>723,1770=>723,1771=>722,1772=>721,1773=>720,1774=>720,1775=>719,1776=>718,1777=>718,1778=>717,1779=>716,1780=>715,1781=>715,1782=>714,1783=>713,1784=>713,1785=>712,1786=>711,1787=>710,1788=>710,1789=>709,1790=>708,1791=>707,1792=>707,1793=>706,1794=>705,1795=>705,1796=>704,1797=>703,1798=>702,1799=>702,1800=>701,1801=>700,1802=>699,1803=>699,1804=>698,1805=>697,1806=>697,1807=>696,1808=>695,1809=>694,1810=>694,1811=>693,1812=>692,1813=>691,1814=>691,1815=>690,1816=>689,1817=>688,1818=>688,1819=>687,1820=>686,1821=>686,1822=>685,1823=>684,1824=>683,1825=>683,1826=>682,1827=>681,1828=>680,1829=>680,1830=>679,1831=>678,1832=>677,1833=>677,1834=>676,1835=>675,1836=>674,1837=>674,1838=>673,1839=>672,1840=>671,1841=>671,1842=>670,1843=>669,1844=>668,1845=>668,1846=>667,1847=>666,1848=>665,1849=>665,1850=>664,1851=>663,1852=>662,1853=>662,1854=>661,1855=>660,1856=>659,1857=>659,1858=>658,1859=>657,1860=>656,1861=>656,1862=>655,1863=>654,1864=>653,1865=>653,1866=>652,1867=>651,1868=>650,1869=>650,1870=>649,1871=>648,1872=>647,1873=>647,1874=>646,1875=>645,1876=>644,1877=>644,1878=>643,1879=>642,1880=>641,1881=>641,1882=>640,1883=>639,1884=>638,1885=>638,1886=>637,1887=>636,1888=>635,1889=>635,1890=>634,1891=>633,1892=>632,1893=>631,1894=>631,1895=>630,1896=>629,1897=>628,1898=>628,1899=>627,1900=>626,1901=>625,1902=>625,1903=>624,1904=>623,1905=>622,1906=>622,1907=>621,1908=>620,1909=>619,1910=>618,1911=>618,1912=>617,1913=>616,1914=>615,1915=>615,1916=>614,1917=>613,1918=>612,1919=>612,1920=>611,1921=>610,1922=>609,1923=>608,1924=>608,1925=>607,1926=>606,1927=>605,1928=>605,1929=>604,1930=>603,1931=>602,1932=>602,1933=>601,1934=>600,1935=>599,1936=>598,1937=>598,1938=>597,1939=>596,1940=>595,1941=>595,1942=>594,1943=>593,1944=>592,1945=>591,1946=>591,1947=>590,1948=>589,1949=>588,1950=>588,1951=>587,1952=>586,1953=>585,1954=>585,1955=>584,1956=>583,1957=>582,1958=>581,1959=>581,1960=>580,1961=>579,1962=>578,1963=>578,1964=>577,1965=>576,1966=>575,1967=>574,1968=>574,1969=>573,1970=>572,1971=>571,1972=>570,1973=>570,1974=>569,1975=>568,1976=>567,1977=>567,1978=>566,1979=>565,1980=>564,1981=>563,1982=>563,1983=>562,1984=>561,1985=>560,1986=>560,1987=>559,1988=>558,1989=>557,1990=>556,1991=>556,1992=>555,1993=>554,1994=>553,1995=>553,1996=>552,1997=>551,1998=>550,1999=>549,2000=>549,2001=>548,2002=>547,2003=>546,2004=>545,2005=>545,2006=>544,2007=>543,2008=>542,2009=>542,2010=>541,2011=>540,2012=>539,2013=>538,2014=>538,2015=>537,2016=>536,2017=>535,2018=>535,2019=>534,2020=>533,2021=>532,2022=>531,2023=>531,2024=>530,2025=>529,2026=>528,2027=>527,2028=>527,2029=>526,2030=>525,2031=>524,2032=>524,2033=>523,2034=>522,2035=>521,2036=>520,2037=>520,2038=>519,2039=>518,2040=>517,2041=>516,2042=>516,2043=>515,2044=>514,2045=>513,2046=>513,2047=>512,2048=>511,2049=>510,2050=>509,2051=>509,2052=>508,2053=>507,2054=>506,2055=>506,2056=>505,2057=>504,2058=>503,2059=>502,2060=>502,2061=>501,2062=>500,2063=>499,2064=>498,2065=>498,2066=>497,2067=>496,2068=>495,2069=>495,2070=>494,2071=>493,2072=>492,2073=>491,2074=>491,2075=>490,2076=>489,2077=>488,2078=>487,2079=>487,2080=>486,2081=>485,2082=>484,2083=>484,2084=>483,2085=>482,2086=>481,2087=>480,2088=>480,2089=>479,2090=>478,2091=>477,2092=>477,2093=>476,2094=>475,2095=>474,2096=>473,2097=>473,2098=>472,2099=>471,2100=>470,2101=>469,2102=>469,2103=>468,2104=>467,2105=>466,2106=>466,2107=>465,2108=>464,2109=>463,2110=>462,2111=>462,2112=>461,2113=>460,2114=>459,2115=>459,2116=>458,2117=>457,2118=>456,2119=>455,2120=>455,2121=>454,2122=>453,2123=>452,2124=>452,2125=>451,2126=>450,2127=>449,2128=>448,2129=>448,2130=>447,2131=>446,2132=>445,2133=>444,2134=>444,2135=>443,2136=>442,2137=>441,2138=>441,2139=>440,2140=>439,2141=>438,2142=>437,2143=>437,2144=>436,2145=>435,2146=>434,2147=>434,2148=>433,2149=>432,2150=>431,2151=>431,2152=>430,2153=>429,2154=>428,2155=>427,2156=>427,2157=>426,2158=>425,2159=>424,2160=>424,2161=>423,2162=>422,2163=>421,2164=>420,2165=>420,2166=>419,2167=>418,2168=>417,2169=>417,2170=>416,2171=>415,2172=>414,2173=>414,2174=>413,2175=>412,2176=>411,2177=>410,2178=>410,2179=>409,2180=>408,2181=>407,2182=>407,2183=>406,2184=>405,2185=>404,2186=>404,2187=>403,2188=>402,2189=>401,2190=>400,2191=>400,2192=>399,2193=>398,2194=>397,2195=>397,2196=>396,2197=>395,2198=>394,2199=>394,2200=>393,2201=>392,2202=>391,2203=>391,2204=>390,2205=>389,2206=>388,2207=>387,2208=>387,2209=>386,2210=>385,2211=>384,2212=>384,2213=>383,2214=>382,2215=>381,2216=>381,2217=>380,2218=>379,2219=>378,2220=>378,2221=>377,2222=>376,2223=>375,2224=>375,2225=>374,2226=>373,2227=>372,2228=>372,2229=>371,2230=>370,2231=>369,2232=>369,2233=>368,2234=>367,2235=>366,2236=>366,2237=>365,2238=>364,2239=>363,2240=>363,2241=>362,2242=>361,2243=>360,2244=>360,2245=>359,2246=>358,2247=>357,2248=>357,2249=>356,2250=>355,2251=>354,2252=>354,2253=>353,2254=>352,2255=>351,2256=>351,2257=>350,2258=>349,2259=>348,2260=>348,2261=>347,2262=>346,2263=>345,2264=>345,2265=>344,2266=>343,2267=>342,2268=>342,2269=>341,2270=>340,2271=>339,2272=>339,2273=>338,2274=>337,2275=>336,2276=>336,2277=>335,2278=>334,2279=>334,2280=>333,2281=>332,2282=>331,2283=>331,2284=>330,2285=>329,2286=>328,2287=>328,2288=>327,2289=>326,2290=>325,2291=>325,2292=>324,2293=>323,2294=>323,2295=>322,2296=>321,2297=>320,2298=>320,2299=>319,2300=>318,2301=>317,2302=>317,2303=>316,2304=>315,2305=>315,2306=>314,2307=>313,2308=>312,2309=>312,2310=>311,2311=>310,2312=>309,2313=>309,2314=>308,2315=>307,2316=>307,2317=>306,2318=>305,2319=>304,2320=>304,2321=>303,2322=>302,2323=>302,2324=>301,2325=>300,2326=>299,2327=>299,2328=>298,2329=>297,2330=>297,2331=>296,2332=>295,2333=>294,2334=>294,2335=>293,2336=>292,2337=>292,2338=>291,2339=>290,2340=>289,2341=>289,2342=>288,2343=>287,2344=>287,2345=>286,2346=>285,2347=>285,2348=>284,2349=>283,2350=>282,2351=>282,2352=>281,2353=>280,2354=>280,2355=>279,2356=>278,2357=>278,2358=>277,2359=>276,2360=>275,2361=>275,2362=>274,2363=>273,2364=>273,2365=>272,2366=>271,2367=>271,2368=>270,2369=>269,2370=>268,2371=>268,2372=>267,2373=>266,2374=>266,2375=>265,2376=>264,2377=>264,2378=>263,2379=>262,2380=>262,2381=>261,2382=>260,2383=>260,2384=>259,2385=>258,2386=>258,2387=>257,2388=>256,2389=>255,2390=>255,2391=>254,2392=>253,2393=>253,2394=>252,2395=>251,2396=>251,2397=>250,2398=>249,2399=>249,2400=>248,2401=>247,2402=>247,2403=>246,2404=>245,2405=>245,2406=>244,2407=>243,2408=>243,2409=>242,2410=>241,2411=>241,2412=>240,2413=>239,2414=>239,2415=>238,2416=>237,2417=>237,2418=>236,2419=>235,2420=>235,2421=>234,2422=>233,2423=>233,2424=>232,2425=>231,2426=>231,2427=>230,2428=>229,2429=>229,2430=>228,2431=>227,2432=>227,2433=>226,2434=>226,2435=>225,2436=>224,2437=>224,2438=>223,2439=>222,2440=>222,2441=>221,2442=>220,2443=>220,2444=>219,2445=>218,2446=>218,2447=>217,2448=>216,2449=>216,2450=>215,2451=>215,2452=>214,2453=>213,2454=>213,2455=>212,2456=>211,2457=>211,2458=>210,2459=>209,2460=>209,2461=>208,2462=>208,2463=>207,2464=>206,2465=>206,2466=>205,2467=>204,2468=>204,2469=>203,2470=>203,2471=>202,2472=>201,2473=>201,2474=>200,2475=>199,2476=>199,2477=>198,2478=>198,2479=>197,2480=>196,2481=>196,2482=>195,2483=>194,2484=>194,2485=>193,2486=>193,2487=>192,2488=>191,2489=>191,2490=>190,2491=>190,2492=>189,2493=>188,2494=>188,2495=>187,2496=>187,2497=>186,2498=>185,2499=>185,2500=>184,2501=>183,2502=>183,2503=>182,2504=>182,2505=>181,2506=>180,2507=>180,2508=>179,2509=>179,2510=>178,2511=>177,2512=>177,2513=>176,2514=>176,2515=>175,2516=>175,2517=>174,2518=>173,2519=>173,2520=>172,2521=>172,2522=>171,2523=>170,2524=>170,2525=>169,2526=>169,2527=>168,2528=>167,2529=>167,2530=>166,2531=>166,2532=>165,2533=>165,2534=>164,2535=>163,2536=>163,2537=>162,2538=>162,2539=>161,2540=>161,2541=>160,2542=>159,2543=>159,2544=>158,2545=>158,2546=>157,2547=>157,2548=>156,2549=>155,2550=>155,2551=>154,2552=>154,2553=>153,2554=>153,2555=>152,2556=>152,2557=>151,2558=>150,2559=>150,2560=>149,2561=>149,2562=>148,2563=>148,2564=>147,2565=>147,2566=>146,2567=>145,2568=>145,2569=>144,2570=>144,2571=>143,2572=>143,2573=>142,2574=>142,2575=>141,2576=>141,2577=>140,2578=>139,2579=>139,2580=>138,2581=>138,2582=>137,2583=>137,2584=>136,2585=>136,2586=>135,2587=>135,2588=>134,2589=>134,2590=>133,2591=>133,2592=>132,2593=>131,2594=>131,2595=>130,2596=>130,2597=>129,2598=>129,2599=>128,2600=>128,2601=>127,2602=>127,2603=>126,2604=>126,2605=>125,2606=>125,2607=>124,2608=>124,2609=>123,2610=>123,2611=>122,2612=>122,2613=>121,2614=>121,2615=>120,2616=>120,2617=>119,2618=>119,2619=>118,2620=>118,2621=>117,2622=>117,2623=>116,2624=>116,2625=>115,2626=>115,2627=>114,2628=>114,2629=>113,2630=>113,2631=>112,2632=>112,2633=>111,2634=>111,2635=>110,2636=>110,2637=>109,2638=>109,2639=>108,2640=>108,2641=>107,2642=>107,2643=>106,2644=>106,2645=>105,2646=>105,2647=>104,2648=>104,2649=>103,2650=>103,2651=>103,2652=>102,2653=>102,2654=>101,2655=>101,2656=>100,2657=>100,2658=>99,2659=>99,2660=>98,2661=>98,2662=>97,2663=>97,2664=>96,2665=>96,2666=>96,2667=>95,2668=>95,2669=>94,2670=>94,2671=>93,2672=>93,2673=>92,2674=>92,2675=>91,2676=>91,2677=>91,2678=>90,2679=>90,2680=>89,2681=>89,2682=>88,2683=>88,2684=>87,2685=>87,2686=>87,2687=>86,2688=>86,2689=>85,2690=>85,2691=>84,2692=>84,2693=>84,2694=>83,2695=>83,2696=>82,2697=>82,2698=>81,2699=>81,2700=>81,2701=>80,2702=>80,2703=>79,2704=>79,2705=>78,2706=>78,2707=>78,2708=>77,2709=>77,2710=>76,2711=>76,2712=>76,2713=>75,2714=>75,2715=>74,2716=>74,2717=>73,2718=>73,2719=>73,2720=>72,2721=>72,2722=>71,2723=>71,2724=>71,2725=>70,2726=>70,2727=>69,2728=>69,2729=>69,2730=>68,2731=>68,2732=>68,2733=>67,2734=>67,2735=>66,2736=>66,2737=>66,2738=>65,2739=>65,2740=>64,2741=>64,2742=>64,2743=>63,2744=>63,2745=>63,2746=>62,2747=>62,2748=>61,2749=>61,2750=>61,2751=>60,2752=>60,2753=>60,2754=>59,2755=>59,2756=>58,2757=>58,2758=>58,2759=>57,2760=>57,2761=>57,2762=>56,2763=>56,2764=>56,2765=>55,2766=>55,2767=>54,2768=>54,2769=>54,2770=>53,2771=>53,2772=>53,2773=>52,2774=>52,2775=>52,2776=>51,2777=>51,2778=>51,2779=>50,2780=>50,2781=>50,2782=>49,2783=>49,2784=>49,2785=>48,2786=>48,2787=>48,2788=>47,2789=>47,2790=>47,2791=>46,2792=>46,2793=>46,2794=>45,2795=>45,2796=>45,2797=>44,2798=>44,2799=>44,2800=>43,2801=>43,2802=>43,2803=>42,2804=>42,2805=>42,2806=>41,2807=>41,2808=>41,2809=>41,2810=>40,2811=>40,2812=>40,2813=>39,2814=>39,2815=>39,2816=>38,2817=>38,2818=>38,2819=>38,2820=>37,2821=>37,2822=>37,2823=>36,2824=>36,2825=>36,2826=>35,2827=>35,2828=>35,2829=>35,2830=>34,2831=>34,2832=>34,2833=>33,2834=>33,2835=>33,2836=>33,2837=>32,2838=>32,2839=>32,2840=>32,2841=>31,2842=>31,2843=>31,2844=>30,2845=>30,2846=>30,2847=>30,2848=>29,2849=>29,2850=>29,2851=>29,2852=>28,2853=>28,2854=>28,2855=>28,2856=>27,2857=>27,2858=>27,2859=>27,2860=>26,2861=>26,2862=>26,2863=>26,2864=>25,2865=>25,2866=>25,2867=>25,2868=>24,2869=>24,2870=>24,2871=>24,2872=>23,2873=>23,2874=>23,2875=>23,2876=>22,2877=>22,2878=>22,2879=>22,2880=>22,2881=>21,2882=>21,2883=>21,2884=>21,2885=>20,2886=>20,2887=>20,2888=>20,2889=>20,2890=>19,2891=>19,2892=>19,2893=>19,2894=>18,2895=>18,2896=>18,2897=>18,2898=>18,2899=>17,2900=>17,2901=>17,2902=>17,2903=>17,2904=>16,2905=>16,2906=>16,2907=>16,2908=>16,2909=>15,2910=>15,2911=>15,2912=>15,2913=>15,2914=>14,2915=>14,2916=>14,2917=>14,2918=>14,2919=>14,2920=>13,2921=>13,2922=>13,2923=>13,2924=>13,2925=>12,2926=>12,2927=>12,2928=>12,2929=>12,2930=>12,2931=>11,2932=>11,2933=>11,2934=>11,2935=>11,2936=>11,2937=>10,2938=>10,2939=>10,2940=>10,2941=>10,2942=>10,2943=>9,2944=>9,2945=>9,2946=>9,2947=>9,2948=>9,2949=>9,2950=>8,2951=>8,2952=>8,2953=>8,2954=>8,2955=>8,2956=>8,2957=>7,2958=>7,2959=>7,2960=>7,2961=>7,2962=>7,2963=>7,2964=>7,2965=>6,2966=>6,2967=>6,2968=>6,2969=>6,2970=>6,2971=>6,2972=>6,2973=>5,2974=>5,2975=>5,2976=>5,2977=>5,2978=>5,2979=>5,2980=>5,2981=>4,2982=>4,2983=>4,2984=>4,2985=>4,2986=>4,2987=>4,2988=>4,2989=>4,2990=>4,2991=>3,2992=>3,2993=>3,2994=>3,2995=>3,2996=>3,2997=>3,2998=>3,2999=>3,3000=>3,3001=>3,3002=>2,3003=>2,3004=>2,3005=>2,3006=>2,3007=>2,3008=>2,3009=>2,3010=>2,3011=>2,3012=>2,3013=>2,3014=>2,3015=>1,3016=>1,3017=>1,3018=>1,3019=>1,3020=>1,3021=>1,3022=>1,3023=>1,3024=>1,3025=>1,3026=>1,3027=>1,3028=>1,3029=>1,3030=>1,3031=>1,3032=>0,3033=>0,3034=>0,3035=>0,3036=>0,3037=>0,3038=>0,3039=>0,3040=>0,3041=>0,3042=>0,3043=>0,3044=>0,3045=>0,3046=>0,3047=>0,3048=>0,3049=>0,3050=>0,3051=>0,3052=>0,3053=>0,3054=>0,3055=>0,3056=>0,3057=>0,3058=>0,3059=>0,3060=>0,3061=>0,3062=>0,3063=>0,3064=>0,3065=>0,3066=>0,3067=>0,3068=>0,3069=>0,3070=>0,3071=>0,3072=>0,3073=>0,3074=>0,3075=>0,3076=>0,3077=>0,3078=>0,3079=>0,3080=>0,3081=>0,3082=>0,3083=>0,3084=>0,3085=>0,3086=>0,3087=>0,3088=>0,3089=>0,3090=>0,3091=>0,3092=>0,3093=>0,3094=>0,3095=>0,3096=>0,3097=>0,3098=>0,3099=>0,3100=>0,3101=>0,3102=>0,3103=>0,3104=>0,3105=>0,3106=>0,3107=>0,3108=>0,3109=>0,3110=>0,3111=>0,3112=>0,3113=>1,3114=>1,3115=>1,3116=>1,3117=>1,3118=>1,3119=>1,3120=>1,3121=>1,3122=>1,3123=>1,3124=>1,3125=>1,3126=>1,3127=>1,3128=>1,3129=>1,3130=>2,3131=>2,3132=>2,3133=>2,3134=>2,3135=>2,3136=>2,3137=>2,3138=>2,3139=>2,3140=>2,3141=>2,3142=>2,3143=>3,3144=>3,3145=>3,3146=>3,3147=>3,3148=>3,3149=>3,3150=>3,3151=>3,3152=>3,3153=>3,3154=>4,3155=>4,3156=>4,3157=>4,3158=>4,3159=>4,3160=>4,3161=>4,3162=>4,3163=>4,3164=>5,3165=>5,3166=>5,3167=>5,3168=>5,3169=>5,3170=>5,3171=>5,3172=>6,3173=>6,3174=>6,3175=>6,3176=>6,3177=>6,3178=>6,3179=>6,3180=>7,3181=>7,3182=>7,3183=>7,3184=>7,3185=>7,3186=>7,3187=>7,3188=>8,3189=>8,3190=>8,3191=>8,3192=>8,3193=>8,3194=>8,3195=>9,3196=>9,3197=>9,3198=>9,3199=>9,3200=>9,3201=>9,3202=>10,3203=>10,3204=>10,3205=>10,3206=>10,3207=>10,3208=>11,3209=>11,3210=>11,3211=>11,3212=>11,3213=>11,3214=>12,3215=>12,3216=>12,3217=>12,3218=>12,3219=>12,3220=>13,3221=>13,3222=>13,3223=>13,3224=>13,3225=>14,3226=>14,3227=>14,3228=>14,3229=>14,3230=>14,3231=>15,3232=>15,3233=>15,3234=>15,3235=>15,3236=>16,3237=>16,3238=>16,3239=>16,3240=>16,3241=>17,3242=>17,3243=>17,3244=>17,3245=>17,3246=>18,3247=>18,3248=>18,3249=>18,3250=>18,3251=>19,3252=>19,3253=>19,3254=>19,3255=>20,3256=>20,3257=>20,3258=>20,3259=>20,3260=>21,3261=>21,3262=>21,3263=>21,3264=>22,3265=>22,3266=>22,3267=>22,3268=>22,3269=>23,3270=>23,3271=>23,3272=>23,3273=>24,3274=>24,3275=>24,3276=>24,3277=>25,3278=>25,3279=>25,3280=>25,3281=>26,3282=>26,3283=>26,3284=>26,3285=>27,3286=>27,3287=>27,3288=>27,3289=>28,3290=>28,3291=>28,3292=>28,3293=>29,3294=>29,3295=>29,3296=>29,3297=>30,3298=>30,3299=>30,3300=>30,3301=>31,3302=>31,3303=>31,3304=>32,3305=>32,3306=>32,3307=>32,3308=>33,3309=>33,3310=>33,3311=>33,3312=>34,3313=>34,3314=>34,3315=>35,3316=>35,3317=>35,3318=>35,3319=>36,3320=>36,3321=>36,3322=>37,3323=>37,3324=>37,3325=>38,3326=>38,3327=>38,3328=>38,3329=>39,3330=>39,3331=>39,3332=>40,3333=>40,3334=>40,3335=>41,3336=>41,3337=>41,3338=>41,3339=>42,3340=>42,3341=>42,3342=>43,3343=>43,3344=>43,3345=>44,3346=>44,3347=>44,3348=>45,3349=>45,3350=>45,3351=>46,3352=>46,3353=>46,3354=>47,3355=>47,3356=>47,3357=>48,3358=>48,3359=>48,3360=>49,3361=>49,3362=>49,3363=>50,3364=>50,3365=>50,3366=>51,3367=>51,3368=>51,3369=>52,3370=>52,3371=>52,3372=>53,3373=>53,3374=>53,3375=>54,3376=>54,3377=>54,3378=>55,3379=>55,3380=>56,3381=>56,3382=>56,3383=>57,3384=>57,3385=>57,3386=>58,3387=>58,3388=>58,3389=>59,3390=>59,3391=>60,3392=>60,3393=>60,3394=>61,3395=>61,3396=>61,3397=>62,3398=>62,3399=>63,3400=>63,3401=>63,3402=>64,3403=>64,3404=>64,3405=>65,3406=>65,3407=>66,3408=>66,3409=>66,3410=>67,3411=>67,3412=>68,3413=>68,3414=>68,3415=>69,3416=>69,3417=>69,3418=>70,3419=>70,3420=>71,3421=>71,3422=>71,3423=>72,3424=>72,3425=>73,3426=>73,3427=>73,3428=>74,3429=>74,3430=>75,3431=>75,3432=>76,3433=>76,3434=>76,3435=>77,3436=>77,3437=>78,3438=>78,3439=>78,3440=>79,3441=>79,3442=>80,3443=>80,3444=>81,3445=>81,3446=>81,3447=>82,3448=>82,3449=>83,3450=>83,3451=>84,3452=>84,3453=>84,3454=>85,3455=>85,3456=>86,3457=>86,3458=>87,3459=>87,3460=>87,3461=>88,3462=>88,3463=>89,3464=>89,3465=>90,3466=>90,3467=>91,3468=>91,3469=>91,3470=>92,3471=>92,3472=>93,3473=>93,3474=>94,3475=>94,3476=>95,3477=>95,3478=>96,3479=>96,3480=>96,3481=>97,3482=>97,3483=>98,3484=>98,3485=>99,3486=>99,3487=>100,3488=>100,3489=>101,3490=>101,3491=>102,3492=>102,3493=>103,3494=>103,3495=>103,3496=>104,3497=>104,3498=>105,3499=>105,3500=>106,3501=>106,3502=>107,3503=>107,3504=>108,3505=>108,3506=>109,3507=>109,3508=>110,3509=>110,3510=>111,3511=>111,3512=>112,3513=>112,3514=>113,3515=>113,3516=>114,3517=>114,3518=>115,3519=>115,3520=>116,3521=>116,3522=>117,3523=>117,3524=>118,3525=>118,3526=>119,3527=>119,3528=>120,3529=>120,3530=>121,3531=>121,3532=>122,3533=>122,3534=>123,3535=>123,3536=>124,3537=>124,3538=>125,3539=>125,3540=>126,3541=>126,3542=>127,3543=>127,3544=>128,3545=>128,3546=>129,3547=>129,3548=>130,3549=>130,3550=>131,3551=>131,3552=>132,3553=>133,3554=>133,3555=>134,3556=>134,3557=>135,3558=>135,3559=>136,3560=>136,3561=>137,3562=>137,3563=>138,3564=>138,3565=>139,3566=>139,3567=>140,3568=>141,3569=>141,3570=>142,3571=>142,3572=>143,3573=>143,3574=>144,3575=>144,3576=>145,3577=>145,3578=>146,3579=>147,3580=>147,3581=>148,3582=>148,3583=>149,3584=>149,3585=>150,3586=>150,3587=>151,3588=>152,3589=>152,3590=>153,3591=>153,3592=>154,3593=>154,3594=>155,3595=>155,3596=>156,3597=>157,3598=>157,3599=>158,3600=>158,3601=>159,3602=>159,3603=>160,3604=>161,3605=>161,3606=>162,3607=>162,3608=>163,3609=>163,3610=>164,3611=>165,3612=>165,3613=>166,3614=>166,3615=>167,3616=>167,3617=>168,3618=>169,3619=>169,3620=>170,3621=>170,3622=>171,3623=>172,3624=>172,3625=>173,3626=>173,3627=>174,3628=>175,3629=>175,3630=>176,3631=>176,3632=>177,3633=>177,3634=>178,3635=>179,3636=>179,3637=>180,3638=>180,3639=>181,3640=>182,3641=>182,3642=>183,3643=>183,3644=>184,3645=>185,3646=>185,3647=>186,3648=>187,3649=>187,3650=>188,3651=>188,3652=>189,3653=>190,3654=>190,3655=>191,3656=>191,3657=>192,3658=>193,3659=>193,3660=>194,3661=>194,3662=>195,3663=>196,3664=>196,3665=>197,3666=>198,3667=>198,3668=>199,3669=>199,3670=>200,3671=>201,3672=>201,3673=>202,3674=>203,3675=>203,3676=>204,3677=>204,3678=>205,3679=>206,3680=>206,3681=>207,3682=>208,3683=>208,3684=>209,3685=>209,3686=>210,3687=>211,3688=>211,3689=>212,3690=>213,3691=>213,3692=>214,3693=>215,3694=>215,3695=>216,3696=>216,3697=>217,3698=>218,3699=>218,3700=>219,3701=>220,3702=>220,3703=>221,3704=>222,3705=>222,3706=>223,3707=>224,3708=>224,3709=>225,3710=>226,3711=>226,3712=>227,3713=>227,3714=>228,3715=>229,3716=>229,3717=>230,3718=>231,3719=>231,3720=>232,3721=>233,3722=>233,3723=>234,3724=>235,3725=>235,3726=>236,3727=>237,3728=>237,3729=>238,3730=>239,3731=>239,3732=>240,3733=>241,3734=>241,3735=>242,3736=>243,3737=>243,3738=>244,3739=>245,3740=>245,3741=>246,3742=>247,3743=>247,3744=>248,3745=>249,3746=>249,3747=>250,3748=>251,3749=>251,3750=>252,3751=>253,3752=>253,3753=>254,3754=>255,3755=>255,3756=>256,3757=>257,3758=>258,3759=>258,3760=>259,3761=>260,3762=>260,3763=>261,3764=>262,3765=>262,3766=>263,3767=>264,3768=>264,3769=>265,3770=>266,3771=>266,3772=>267,3773=>268,3774=>268,3775=>269,3776=>270,3777=>271,3778=>271,3779=>272,3780=>273,3781=>273,3782=>274,3783=>275,3784=>275,3785=>276,3786=>277,3787=>278,3788=>278,3789=>279,3790=>280,3791=>280,3792=>281,3793=>282,3794=>282,3795=>283,3796=>284,3797=>285,3798=>285,3799=>286,3800=>287,3801=>287,3802=>288,3803=>289,3804=>289,3805=>290,3806=>291,3807=>292,3808=>292,3809=>293,3810=>294,3811=>294,3812=>295,3813=>296,3814=>297,3815=>297,3816=>298,3817=>299,3818=>299,3819=>300,3820=>301,3821=>302,3822=>302,3823=>303,3824=>304,3825=>304,3826=>305,3827=>306,3828=>307,3829=>307,3830=>308,3831=>309,3832=>309,3833=>310,3834=>311,3835=>312,3836=>312,3837=>313,3838=>314,3839=>315,3840=>315,3841=>316,3842=>317,3843=>317,3844=>318,3845=>319,3846=>320,3847=>320,3848=>321,3849=>322,3850=>323,3851=>323,3852=>324,3853=>325,3854=>325,3855=>326,3856=>327,3857=>328,3858=>328,3859=>329,3860=>330,3861=>331,3862=>331,3863=>332,3864=>333,3865=>334,3866=>334,3867=>335,3868=>336,3869=>336,3870=>337,3871=>338,3872=>339,3873=>339,3874=>340,3875=>341,3876=>342,3877=>342,3878=>343,3879=>344,3880=>345,3881=>345,3882=>346,3883=>347,3884=>348,3885=>348,3886=>349,3887=>350,3888=>351,3889=>351,3890=>352,3891=>353,3892=>354,3893=>354,3894=>355,3895=>356,3896=>357,3897=>357,3898=>358,3899=>359,3900=>360,3901=>360,3902=>361,3903=>362,3904=>363,3905=>363,3906=>364,3907=>365,3908=>366,3909=>366,3910=>367,3911=>368,3912=>369,3913=>369,3914=>370,3915=>371,3916=>372,3917=>372,3918=>373,3919=>374,3920=>375,3921=>375,3922=>376,3923=>377,3924=>378,3925=>378,3926=>379,3927=>380,3928=>381,3929=>381,3930=>382,3931=>383,3932=>384,3933=>384,3934=>385,3935=>386,3936=>387,3937=>387,3938=>388,3939=>389,3940=>390,3941=>391,3942=>391,3943=>392,3944=>393,3945=>394,3946=>394,3947=>395,3948=>396,3949=>397,3950=>397,3951=>398,3952=>399,3953=>400,3954=>400,3955=>401,3956=>402,3957=>403,3958=>404,3959=>404,3960=>405,3961=>406,3962=>407,3963=>407,3964=>408,3965=>409,3966=>410,3967=>410,3968=>411,3969=>412,3970=>413,3971=>414,3972=>414,3973=>415,3974=>416,3975=>417,3976=>417,3977=>418,3978=>419,3979=>420,3980=>420,3981=>421,3982=>422,3983=>423,3984=>424,3985=>424,3986=>425,3987=>426,3988=>427,3989=>427,3990=>428,3991=>429,3992=>430,3993=>431,3994=>431,3995=>432,3996=>433,3997=>434,3998=>434,3999=>435,4000=>436,4001=>437,4002=>437,4003=>438,4004=>439,4005=>440,4006=>441,4007=>441,4008=>442,4009=>443,4010=>444,4011=>444,4012=>445,4013=>446,4014=>447,4015=>448,4016=>448,4017=>449,4018=>450,4019=>451,4020=>452,4021=>452,4022=>453,4023=>454,4024=>455,4025=>455,4026=>456,4027=>457,4028=>458,4029=>459,4030=>459,4031=>460,4032=>461,4033=>462,4034=>462,4035=>463,4036=>464,4037=>465,4038=>466,4039=>466,4040=>467,4041=>468,4042=>469,4043=>469,4044=>470,4045=>471,4046=>472,4047=>473,4048=>473,4049=>474,4050=>475,4051=>476,4052=>477,4053=>477,4054=>478,4055=>479,4056=>480,4057=>480,4058=>481,4059=>482,4060=>483,4061=>484,4062=>484,4063=>485,4064=>486,4065=>487,4066=>487,4067=>488,4068=>489,4069=>490,4070=>491,4071=>491,4072=>492,4073=>493,4074=>494,4075=>495,4076=>495,4077=>496,4078=>497,4079=>498,4080=>498,4081=>499,4082=>500,4083=>501,4084=>502,4085=>502,4086=>503,4087=>504,4088=>505,4089=>506,4090=>506,4091=>507,4092=>508,4093=>509,4094=>509,4095=>510);
signal coef : integer range 0 to 1023;		-- Koeffizient der Funktion aus Koeffiziententabelle
signal c : integer range 0 to 1023 := 0;	-- Z�hler des Taktteilers f�r f_ref
signal pwm_counter : integer := 0;			-- z�hlt wie viel Takte in aktueller Periode vergangen sind

begin
-- Generierung der Referenzfrequenz mit 48.828 kHz
f_ref_generierung: process
begin
	-- jeden 1023ten Takt f_ref für einen Takt auf high -> f_ref mit 50 MHz / 1023 = 48.828 kHz
	if (c = 1023) then
		c <= 0;
		f_ref <= '1';
	else
		c <= c + 1;
		f_ref <= '0';
	end if;

	wait for 20 ns;
end process f_ref_generierung;

-- Generierung des Phasenwerts
phasenakkumulator: process(f_ref)
begin
	-- addiert einmal pro Periode von f_ref f_sel zur Phase
	if rising_edge(f_ref) then
		if (phase + f_sel < 4096) then
			phase <= phase + f_sel;
		else
			phase <= phase + f_sel - 4096;
		end if;
	end if;
end process phasenakkumulator;

-- Generierung des PWM-Signals aus Koeffizienten
pwm_generierung: process
begin
	-- neue Periode beginnt wenn f_ref auslöst -> Zähler zurücksetzen
	if (pwm_counter >= 1023) then
		pwm_counter <= 0;
		coef <= coef_table(phase);
	else
		pwm_counter <= pwm_counter + 1;
	end if;
	-- die ersten coef Takte ist der PWM-Ausgang auf high, danach auf low
	if (pwm_counter <= coef) then
		pwm_out <= '1';
	else
		pwm_out <= '0';
	end if;

	wait for 20 ns;
end process pwm_generierung;

end algorithmisch;