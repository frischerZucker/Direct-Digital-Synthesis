library ieee;

package coef_table_package is
	type coef_table_t is array (0 to 4095) of integer;
end coef_table_package;

package body coef_table_package is

end coef_table_package;